////////////////////////////////////////////////////////////////////////
// Developer Name : Mohsan Naeem 
// Contact info   : mohsannaeem1576@gmail.com
// Module Name    : ahb_env_pkg
// Description    : Dummy env_pkg which can be used to create new env_pkg
///////////////////////////////////////////////////////////////////////
package ahb_env_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"
    import ahb_seq_pkg::*;
   `include "ahb_mst_agent_config.sv"
   `include "ahb_slv_agent_config.sv"
   `include "ahb_env_config.sv"
   `include "ahb_mst_sequencer.sv"
   `include "ahb_mst_driver.sv"
   `include "ahb_mst_agent.sv"
   `include "ahb_slv_sequencer.sv"
   `include "ahb_slv_driver.sv"
   `include "ahb_slv_agent.sv"
   `include "ahb_env.sv"
endpackage