////////////////////////////////////////////////////////////////////////
// Developer Name : Mohsan Naeem 
// Contact info   : mohsannaeem1576@gmail.com
// Module Name    : ahb_seq_pkg
// Description    : Dummy seq_pkg which can be used to create new seq_pkg
///////////////////////////////////////////////////////////////////////
package ahb_seq_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "ahb_mst_seq_item.sv"
	`include "ahb_mst_base_sequence.sv"
  `include "ahb_slv_seq_item.sv"
  `include "ahb_slv_base_sequence.sv"
endpackage