////////////////////////////////////////////////////////////////////////
// Developer Name : Mohsan Naeem 
// Contact info   : mohsannaeem1576@gmail.com
// Module Name    : ahb_test_pkg
// Description    : Dummy Test Package which can be used to create new test pkg
///////////////////////////////////////////////////////////////////////
package ahb_test_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import ahb_seq_pkg::*;
    import ahb_env_pkg::*;
    `include "ahb_base_test.sv"
endpackage